module adder(a0,a1,a2,a3,sum);
input[7:0] a0,a1,a2,a3,sum;
reg[7:0] sum;
and()
endmodule