module adder(a0,a1,a2,a3,cout,sum);
input[7:0] a0,a1,a2,a3;
output[1:0] cout;
output[7:0] sum;
reg[7:0] sum;
reg c0,c1,c2;
reg[1:0] cout;
reg[7:0] tmp0,tmp1;
always@(a0 or a1 or a2 or a3)
begin
	{c0,tmp0} = a0+a1;
	{c1,tmp1} = a2+tmp0;
	{c2,sum} = tmp1+a3;
	cout = c2+c0+c1;
end
endmodule